`timescale 1ns/10ps

/* resource counter for nor gates
 */

module global_vars;
initial
integer count=0;
endmodule
