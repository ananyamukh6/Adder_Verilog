`timescale 1ns/10ps

/* resource counter for nor gates
 */

module global_vars;
integer count;
initial
count=0;
endmodule
